// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Apr  2023  
// (c) Technion IIT, Department of Electrical Engineering 2023 

module	ShieldMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic collision, //changed random_hart to collision
					input logic startOfFrame,				
					input monster_barrier_collision,
			
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */


// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 16*16 and use only the top left 16*15 squares 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the  understanding 
int flag = 0;

logic [0:63] [0:63] [3:0]  MazeBitMapMask ;  //matrix the each 1,2,0 represents a diffrent bitmap from bellow

logic [0:63] [0:63] [3:0]  MazeDefaultBitMapMask= // defult table to load on reset 
{{128'h00000000000000000000000000000000},     
 {128'h00000000000000000000000000000000},
 {128'h00000000110000000001100000000000},
 {128'h00000000000000000000000000000000},
 {128'h00110000000000000000000000000000},
 {128'h00000000000000000110000000000000},
 {128'h00000001100000000000000000000000},
 {128'h00000000000000000000000011000000},
 {128'h00000000000000000000000000000000},
 {128'h00000000000000000000000000000000},
 {128'h00110011011001100000000000000000},
 {128'h00000000000000000000000000110000},
 {128'h00000000000000000000000000000000},
 {128'h00000000000001100000000000000000},
 {128'h00000000000000000000000000000000},
 {128'h00000000000000000000000000000000}};


 
 
//first is before second is after collision
 logic [1:0] [0:15] [0:15] [7:0]  object_colors  = {
{{8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h00,8'h24,8'h24,8'h00,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00},
	{8'h00,8'h24,8'h1a,8'hbf,8'h3e,8'hbf,8'h24,8'hdf,8'hb6,8'h24,8'hbf,8'h3e,8'hbf,8'h1a,8'h24,8'h00},
	{8'h24,8'h1a,8'hb6,8'hba,8'hff,8'hb6,8'h24,8'hb6,8'hdf,8'h24,8'hb6,8'hdf,8'hb6,8'h3e,8'h1a,8'h24},
	{8'h24,8'hbf,8'hdf,8'h3e,8'h1a,8'h3e,8'h24,8'hba,8'hb6,8'h24,8'h1a,8'h1a,8'h3e,8'hbf,8'hbf,8'h24},
	{8'h24,8'hbf,8'hbf,8'h3e,8'hbf,8'h1a,8'h24,8'hdf,8'hba,8'h24,8'h1a,8'hbf,8'h1a,8'hdf,8'h3e,8'h24},
	{8'h24,8'hbf,8'hb6,8'h3e,8'h1a,8'hb6,8'h24,8'hba,8'hb6,8'h24,8'hb6,8'h1a,8'hbf,8'hba,8'hbf,8'h24},
	{8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h1a,8'h24,8'h24,8'hbf,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00},
	{8'h24,8'hb6,8'hba,8'hdf,8'hb6,8'hba,8'h24,8'h1a,8'hbf,8'h24,8'hb6,8'hdf,8'hba,8'hb6,8'hb6,8'h24},
	{8'h24,8'hba,8'hdf,8'hb6,8'hba,8'hdf,8'h24,8'hbf,8'h3e,8'h24,8'hdf,8'hb6,8'hb6,8'hba,8'hdf,8'h24},
	{8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h3e,8'h24,8'h24,8'hbf,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00},
	{8'h24,8'hff,8'hb6,8'h3e,8'h1a,8'hb6,8'h24,8'hdf,8'hb6,8'h24,8'hb6,8'h1a,8'h3e,8'hdf,8'hbf,8'h24},
	{8'h24,8'hbf,8'h1a,8'hbf,8'h3e,8'h1a,8'h24,8'hb6,8'hba,8'h24,8'h1a,8'h1a,8'hbf,8'hb6,8'h3e,8'h24},
	{8'h24,8'hbf,8'hdf,8'h3e,8'h1a,8'h3e,8'h24,8'hba,8'hdf,8'h24,8'h1a,8'hff,8'h1a,8'hbf,8'hbf,8'h24},
	{8'h24,8'h1a,8'hba,8'hdf,8'hbf,8'hb6,8'h24,8'hdf,8'hb6,8'h24,8'hb6,8'hdf,8'hdf,8'hba,8'h1a,8'h24},
	{8'h00,8'h24,8'h1a,8'hbf,8'h3e,8'hbf,8'h24,8'hb6,8'hdf,8'h24,8'hbf,8'h3e,8'hbf,8'h1a,8'h24,8'h00},
	{8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h00,8'h24,8'h24,8'h00,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00}
	},
	
{{8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00},
	{8'h00,8'h24,8'h1a,8'hbf,8'h3e,8'hbf,8'hbf,8'h3e,8'hbf,8'hbf,8'hbf,8'h3e,8'hbf,8'h1a,8'h24,8'h00},
	{8'h24,8'h1a,8'hb6,8'hba,8'hdf,8'hff,8'h3e,8'hba,8'hba,8'hdf,8'hbf,8'hdf,8'hb6,8'hdf,8'h1a,8'h24},
	{8'h24,8'hbf,8'hdf,8'h3e,8'h1a,8'h3e,8'h1a,8'h1a,8'hbf,8'h3e,8'h1a,8'h1a,8'h3e,8'hbf,8'hbf,8'h24},
	{8'h24,8'hbf,8'hbf,8'hff,8'hbf,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'hbf,8'h1a,8'hdf,8'h3e,8'h24},
	{8'h24,8'hbf,8'h1a,8'h3e,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hbf,8'hba,8'hbf,8'h24},
	{8'h24,8'h3e,8'hdf,8'h1a,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h3e,8'hb6,8'hbf,8'h24},
	{8'h24,8'hbf,8'hba,8'h3e,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hbf,8'hdf,8'hbf,8'h24},
	{8'h24,8'hbf,8'hb6,8'hbf,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h1a,8'hba,8'h3e,8'h24},
	{8'h24,8'h3e,8'hdf,8'h1a,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h1a,8'hbf,8'hbf,8'h24},
	{8'h24,8'hbf,8'hbf,8'h3e,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h3e,8'hdf,8'hbf,8'h24},
	{8'h24,8'hbf,8'hb6,8'hbf,8'h3e,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h1a,8'hbf,8'hb6,8'h3e,8'h24},
	{8'h24,8'hbf,8'hdf,8'h3e,8'h1a,8'h3e,8'h1a,8'hbf,8'h1a,8'h3e,8'h1a,8'h3e,8'h1a,8'hbf,8'hbf,8'h24},
	{8'h24,8'h1a,8'hba,8'hdf,8'hbf,8'hff,8'hdf,8'hba,8'hb6,8'hdf,8'hbf,8'hdf,8'hdf,8'hba,8'h1a,8'h24},
	{8'h00,8'h24,8'h1a,8'hbf,8'h3e,8'hbf,8'h3e,8'hbf,8'hbf,8'h3e,8'hbf,8'h3e,8'hbf,8'h1a,8'h24,8'h00},
	{8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00}}
	};
 

typedef enum logic [1:0] {
    COL_ST,           // collision
    PROCESSING_ST // startOfFrame activity-after all data collected 
} state_t;
state_t SM_Shield;

always_ff @(posedge clk or negedge resetN) begin : fsm_sync_proc
    if (resetN == 1'b0) begin 
        SM_Shield <= COL_ST; 
        RGBout <=	8'h00;
		  MazeBitMapMask  <=  MazeDefaultBitMapMask ;  //  copy default tabel 
		  flag <= 0;    
    end else begin
     RGBout <= TRANSPARENT_ENCODING ; // default 
        case (SM_Shield)
            //------------
            COL_ST: begin // position interpolate 
                if (collision == 1'b1 && MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'h1 && flag == 0) begin	//first hit					
						MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h2;
						flag <= 1;	
						SM_Shield <= PROCESSING_ST;	
						end			 
				 else if (collision == 1'b1 && MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'h2 && flag == 0) begin //second hit
						MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h0;
						flag <= 1;
						SM_Shield <= PROCESSING_ST;
						end				  					
            end
        
            //------------------------
            PROCESSING_ST: begin // state to proccess information
                
					 if(startOfFrame) begin
					 SM_Shield <= COL_ST; 
					 flag <= !flag;
					 end
				end
        endcase // case 
    
						if (InsideRectangle == 1'b1 )	
						begin 
							case (MazeBitMapMask[offsetY[8:5]][offsetX[8:5]])
								 4'h0 : RGBout <= TRANSPARENT_ENCODING ; //transperent
								 4'h1 : RGBout <= object_colors[!collision][offsetY[4:0]][offsetX[4:0]]; //shield full hp
								 4'h2 : RGBout <= object_colors[collision][offsetY[4:0]][offsetX[4:0]] ; //shield half hp
								 default:  RGBout <= TRANSPARENT_ENCODING ; 
							endcase						
						end 
					end
end // end fsm_sync
//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule



