//
// coding convention dudy December 2018
// (c) Technion IIT, Department of Electrical Engineering 2021
// generating a number bitmap 



module NumbersBitMapSecond	(	
					input		logic	clk,
					input		logic	resetN,
			    	input 	logic	[10:0] offsetX,// offset from top left  position 
					input 	logic	[10:0] offsetY,
					input 	logic got_hit,
					input 	logic startOfFrame,
					output	logic				drawingRequest,	    								 
					output	logic	[7:0]		RGBout
);
// generating a smily bitmap 
parameter  logic	[7:0] digit_color = 8'hff ; //set the color of the digit 
int hp =100;
bit [0:4] [0:31] [0:63] hp_bitmap  = {



{64'b	0000000011100000000000111110000000000000111110000000000000000000,
 64'b	0000000111100000000011111111100000000011111111100000000000000000,
 64'b	0000011111100000000011111111100000000011111111100000000000000000,
 64'b	0000111111100000000111111111110000000111111111110000000000000000,
 64'b	0001111111100000001111100111110000001111100111110000000000000000,
 64'b	0011111111100000001110000011111000001110000011111000000000000000,
 64'b	0111111011100000011110000001111000011110000001111000000000000000,
 64'b	0111100011100000011110000001111000011110000001111000000000000000,
 64'b	0111000011100000111110000001111100111110000001111100000000000000,
 64'b	0010000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000000111100111100000000111100000000000000,
 64'b	0000000011100000111100000001111000111100000001111000000000000000,
 64'b	0000000011100000111110000001111000111110000001111000000000000000,
 64'b	0000000011100000011111000011111000011111000011111000000000000000,
 64'b	0000000011100000011111000011110000011111000011110000000000000000,
 64'b	0000000011100000001111100111110000001111100111110000000000000000,
 64'b	0111111111111111001111111111100000001111111111100000000000000000,
 64'b	0111111111111111000111111111100000000111111111100000000000000000,
 64'b	0111111111111111000011111111000000000011111111000000000000000000,
 64'b	0111111111111111000001111100000000000001111100000000000000000000,
},


{64'b	0000000000000000111111111111111100011111111111111100000000000000,
 64'b	0000000000000000111111111111111100011111111111111100000000000000,
 64'b	0000000000000000111111111111111100011111111111111000000000000000,
 64'b	0000000000000000111111111111111100011111111111110000000000000000,
 64'b	0000000000000000110000000000111100011110000000000000000000000000,
 64'b	0000000000000000100000000001111100011110000000000000000000000000,
 64'b	0000000000000000000000000001111100011110000000000000000000000000,
 64'b	0000000000000000000000000001111000011110000000000000000000000000,
 64'b	0000000000000000000000000011111000011110000000000000000000000000,
 64'b	0000000000000000000000000011110000011110000000000000000000000000,
 64'b	0000000000000000000000000111110000011110000000000000000000000000,
 64'b	0000000000000000000000000111100000011111111110000000000000000000,
 64'b	0000000000000000000000001111100000011111111111100000000000000000,
 64'b	0000000000000000000000001111100000011111111111100000000000000000,
 64'b	0000000000000000000000001111100000011111111111110000000000000000,
 64'b	0000000000000000000000001111100000001111111111111000000000000000,
 64'b	0000000000000000000000001111000000000000000111111000000000000000,
 64'b	0000000000000000000000001111000000000000000011111100000000000000,
 64'b	0000000000000000000000001110000000000000000001111100000000000000,
 64'b	0000000000000000000000001110000000000000000001111100000000000000,
 64'b	0000000000000000000000011110000000000000000000111100000000000000,
 64'b	0000000000000000000000011110000000000000000000111100000000000000,
 64'b	0000000000000000000000111100000000000000000000111100000000000000,
 64'b	0000000000000000000000111100000000000000000001111100000000000000,
 64'b	0000000000000000000001111000000000000000000001111100000000000000,
 64'b	0000000000000000000001111000000000100000000011111000000000000000,
 64'b	0000000000000000000011111000000000110000000111111000000000000000,
 64'b	0000000000000000000011110000000000111110001111110000000000000000,
 64'b	0000000000000000000011110000000000111111111111100000000000000000,
 64'b	0000000000000000000111110000000000111111111111100000000000000000,
 64'b	0000000000000000000111110000000000111111111111000000000000000000,
 64'b	0000000000000000000111110000000000000111111100000000000000000000,
},

{64'b	0000000000000000000111111111111111000000001111100000000000000000,
 64'b	0000000000000000000111111111111111000000111111111000000000000000,
 64'b	0000000000000000000111111111111110000000111111111000000000000000,
 64'b	0000000000000000000111111111111100000001111111111100000000000000,
 64'b	0000000000000000000111100000000000000011111001111100000000000000,
 64'b	0000000000000000000111100000000000000011100000111110000000000000,
 64'b	0000000000000000000111100000000000000111100000011110000000000000,
 64'b	0000000000000000000111100000000000000111100000011110000000000000,
 64'b	0000000000000000000111100000000000001111100000011111000000000000,
 64'b	0000000000000000000111100000000000001111000000001111000000000000,
 64'b	0000000000000000000111100000000000001111000000001111000000000000,
 64'b	0000000000000000000111111111100000001111000000001111000000000000,
 64'b	0000000000000000000111111111111000001111000000001111000000000000,
 64'b	0000000000000000000111111111111000001111000000001111000000000000,
 64'b	0000000000000000000111111111111100001111000000001111000000000000,
 64'b	0000000000000000000011111111111110001111000000001111000000000000,
 64'b	0000000000000000000000000001111110001111000000001111000000000000,
 64'b	0000000000000000000000000000111111001111000000001111000000000000,
 64'b	0000000000000000000000000000011111001111000000001111000000000000,
 64'b	0000000000000000000000000000011111001111000000001111000000000000,
 64'b	0000000000000000000000000000001111001111000000001111000000000000,
 64'b	0000000000000000000000000000001111001111000000001111000000000000,
 64'b	0000000000000000000000000000001111001111000000001111000000000000,
 64'b	0000000000000000000000000000011111001111000000011110000000000000,
 64'b	0000000000000000000000000000011111001111100000011110000000000000,
 64'b	0000000000000000001000000000111110000111110000111110000000000000,
 64'b	0000000000000000001100000001111110000111110000111100000000000000,
 64'b	0000000000000000001111100011111100000011111001111100000000000000,
 64'b	0000000000000000001111111111111000000011111111111000000000000000,
 64'b	0000000000000000001111111111111000000001111111111000000000000000,
 64'b	0000000000000000001111111111110000000000111111110000000000000000,
 64'b	0000000000000000000001111111000000000000011111000000000000000000,
},

{64'b	0000000000000000000001111111000000001111111111111110000000000000,
 64'b	0000000000000000000011111111100000001111111111111110000000000000,
 64'b	0000000000000000001111111111110000001111111111111100000000000000,
 64'b	0000000000000000011111111111110000001111111111111000000000000000,
 64'b	0000000000000000011111100111111000001111000000000000000000000000,
 64'b	0000000000000000011110000111111000001111000000000000000000000000,
 64'b	0000000000000000011100000011111100001111000000000000000000000000,
 64'b	0000000000000000000000000001111100001111000000000000000000000000,
 64'b	0000000000000000000000000001111100001111000000000000000000000000,
 64'b	0000000000000000000000000001111100001111000000000000000000000000,
 64'b	0000000000000000000000000001111000001111000000000000000000000000,
 64'b	0000000000000000000000000011111000001111111111000000000000000000,
 64'b	0000000000000000000000000011111000001111111111110000000000000000,
 64'b	0000000000000000000000000011110000001111111111110000000000000000,
 64'b	0000000000000000000000000111110000001111111111111000000000000000,
 64'b	0000000000000000000000000111110000000111111111111100000000000000,
 64'b	0000000000000000000000000111110000000000000011111100000000000000,
 64'b	0000000000000000000000000111100000000000000001111110000000000000,
 64'b	0000000000000000000000000111000000000000000000111110000000000000,
 64'b	0000000000000000000000001110000000000000000000111110000000000000,
 64'b	0000000000000000000000011110000000000000000000011110000000000000,
 64'b	0000000000000000000000111100000000000000000000011110000000000000,
 64'b	0000000000000000000001111000000000000000000000011110000000000000,
 64'b	0000000000000000000011111000000000000000000000111110000000000000,
 64'b	0000000000000000000011111000000000000000000000111110000000000000,
 64'b	0000000000000000000111110000000000010000000001111100000000000000,
 64'b	0000000000000000001111100000000010011000000011111100000000000000,
 64'b	0000000000000000011111000000000110011111000111111000000000000000,
 64'b	0000000000000000011111111111111110011111111111110000000000000000,
 64'b	0000000000000000011111111111111110011111111111110000000000000000,
 64'b	0000000000000000011111111111111110011111111111100000000000000000,
 64'b	0000000000000000011111111111111110000011111110000000000000000000,
},
{64'b	0000000000000000000000001111100000000000001111100000000000000000,
 64'b	0000000000000000000000111111111000000000111111111000000000000000,
 64'b	0000000000000000000000111111111000000000111111111000000000000000,
 64'b 0000000000000000000001111111111100000001111111111100000000000000,
 64'b 0000000000000000000011111001111100000011111001111100000000000000,
 64'b 0000000000000000000011100000111110000011100000111110000000000000,
 64'b 0000000000000000000111100000011110000111100000011110000000000000,
 64'b 0000000000000000000111100000011110000111100000011110000000000000,
 64'b 0000000000000000001111100000011111100111100000011111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000001111001111000000001111000000000000,
 64'b 0000000000000000001111000000011110001111000000011110000000000000,
 64'b 0000000000000000001111100000011110001111100000011110000000000000,
 64'b 0000000000000000000111110000111110000111110000111110000000000000,
 64'b 0000000000000000000111110000111100000111110000111100000000000000,
 64'b 0000000000000000000011111001111100000011111001111100000000000000,
 64'b 0000000000000000000011111111111000000011111111111000000000000000,
 64'b 0000000000000000000001111111111000000001111111111000000000000000,
 64'b 0000000000000000000000111111110000000000111111110000000000000000,
 64'b 0000000000000000000000011111000000000000011111000000000000000000,

}};

typedef enum logic [1:0] {
    COL_ST,           // collision
    PROCESSING_ST // startOfFrame activity-after all data collected 
} state_t;
state_t SM_HP;

always_ff @(posedge clk or negedge resetN) begin : fsm_sync_proc
    if (resetN == 1'b0) begin 
        drawingRequest <= (hp_bitmap[0][offsetY][offsetX]);
		  SM_HP <= COL_ST;    
    end else begin     
        case (SM_HP)
            //------------
            COL_ST: begin // position interpolate 
                if (got_hit && hp == 100) begin	//first hit					
						hp <= 75;
						SM_HP <= PROCESSING_ST;	
						end			 
				 else if (got_hit && hp == 75) begin //second hit
						hp <= 50;
						SM_HP <= PROCESSING_ST;
						end
				 else if (got_hit  && hp == 50) begin //second hit
						hp <= 25;
						SM_HP <= PROCESSING_ST;
						end
				  	else if (got_hit  && hp == 25) begin //second hit
						hp <= 0;
						SM_HP <= PROCESSING_ST;
						end		
            end
        
            //------------------------
            PROCESSING_ST: begin // state to proccess information
                
					 if(startOfFrame) begin
					 SM_HP <= COL_ST; 
					 end
				end
        endcase // case   
							case (hp)
								 100 : drawingRequest <= (hp_bitmap[0][offsetY][offsetX]); //full hp
								 75 : drawingRequest <= (hp_bitmap[1][offsetY][offsetX]); //75hp
								 50 : drawingRequest <= (hp_bitmap[2][offsetY][offsetX]); //50
								 25 : drawingRequest <= (hp_bitmap[3][offsetY][offsetX]); //25
								 0 : drawingRequest <= (hp_bitmap[4][offsetY][offsetX]); //00
								 
								 default:  drawingRequest <= (hp_bitmap[0][offsetY][offsetX]); 
							endcase						
						
					end
end // end fsm_sync
//==----------------------------------------------------------------------------------------------------------------=
  

assign RGBout = digit_color ; // this is a fixed color 

endmodule