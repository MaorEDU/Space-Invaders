{
16'b 1110000000000111,
16'b 1110000000000111, 
16'b 1110000000000111,
16'b 1110000000000111,
16'b 1110000000000111,
16'b 1110000000000111,
16'b 1111111111111111,
16'b 1111111111111111,
16'b 1110000000000111,
16'b 1110000000000111,
16'b 1110000000000111,
16'b 1110000000000111,
16'b 1110000000000111,
16'b 1110000000000111,
16'b 1110000000000111,
16'b 1110000000000111
},
	
{
16'b 1111111111111111,
16'b 1111111111111111,
16'b 1110000000000011,
16'b 1110000000000011,
16'b 1110000000000011,
16'b 1110000000000011,
16'b 1111111111111111,
16'b 1111111111111111, 
16'b 1110000000000000,
16'b 1110000000000000,
16'b 1110000000000000,
16'b 1110000000000000,
16'b 1110000000000000,
16'b 1110000000000000,
16'b 1110000000000000,
16'b 1110000000000000
},
 
 {
16'b 0000000000000000,
16'b 0000000000000000,
16'b 0000000000000000,
16'b 0000000000000000, 
16'b 0000000000000000,
16'b 0000011100000000,
16'b 0000011100000000,
16'b 0000011100000000,
16'b 0000011100000000,
16'b 0000000000000000,
16'b 0000000000000000,
16'b 0000011100000000,
16'b 0000011100000000,
16'b 0000011100000000,
16'b 0000011100000000,
16'b 0000000000000000
}};