//
// coding convention dudy December 2018
// (c) Technion IIT, Department of Electrical Engineering 2021
// generating a number bitmap 



module NumbersBitMap	(	
					input		logic	clk,
					input		logic	resetN,
			    	input 	logic	[10:0] offsetX,// offset from top left  position 
					input 	logic	[10:0] offsetY,

					output	logic				drawingRequest,	    								 
					output	logic	[7:0]		RGBout
);
// generating a smily bitmap 
parameter  logic	[7:0] digit_color = 8'hff ; //set the color of the digit 

bit [0:31] [0:63] hp_bitmap  = {



{64'b 00000000011110000000011110001111111111111110000000000000000000,
 64'b 00000000011110000000011110001111111111111110000000000000000000,
 64'b 00000000011110000000011110001111111111111110000000000000000000,
 64'b 00000000011110000000011110001111111111111110000000000000000000,
 64'b 00000000011110000000011110001111100000011110000000000000000000,
 64'b 00000000011110000000011110001111000000001110000000000000000000,
 64'b 00000000011110000000011110001111000000001110000000000000000000,
 64'b 00000000011110000000011110001111000000001110000000000000000000,
 64'b 00000000011110000000011110001111000000001110000000000000000000,
 64'b 00000000011110000000011110001111000000001110000000001100000000,
 64'b 00000000011110000000011110001111000000001110000000011110000000,
 64'b 00000000011110000000011110001111100000011110000000111111000000,
 64'b 00000000011110000000011110001111111111111100000000111111000000,
 64'b 00000000011110000000011110001111111111111100000000011110000000,
 64'b 00000000011110000000011110001111111111111000000000001100000000,
 64'b 00000000011111111111111110001111000000000000000000000000000000,
 64'b 00000000011111111111111110001111000000000000000000000000000000,
 64'b 00000000011111111111111110001111000000000000000000000000000000,
 64'b 00000000011111111111111110001111000000000000000000001100000000,
 64'b 00000000011110000000011110001111000000000000000000011110000000,
 64'b 00000000011110000000011110001111000000000000000000111111000000,
 64'b 00000000011110000000011110001111000000000000000000111111000000,
 64'b 00000000011110000000011110001111000000000000000000011110000000,
 64'b 00000000011110000000011110001111000000000000000000001100000000,
 64'b 00000000011110000000011110001111000000000000000000000000000000,
 64'b 00000000011110000000011110001111000000000000000000000000000000,
 64'b 00000000011110000000011110001111000000000000000000000000000000,
 64'b 00000000011110000000011110001111000000000000000000000000000000,
 64'b 00000000011110000000011110001111000000000000000000000000000000,
 64'b 00000000011110000000011110001111000000000000000000000000000000,
 64'b 00000000011110000000011110001111000000000000000000000000000000,
 64'b 00000000011110000000011110001111000000000000000000000000000000,
}};



// pipeline (ff) to get the pixel color from the array 	 
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
			drawingRequest <= (hp_bitmap[offsetY][offsetX]);
	end
	else 
		drawingRequest <= (hp_bitmap[offsetY][offsetX]);

end


assign RGBout = digit_color ; // this is a fixed color 

endmodule